LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY MAQUINA_DE_ESTADOS IS
	PORT (botao,clk: IN  STD_LOGIC;
          saida:BUFFER STD_LOGIC);
END ENTITY;
    
ARCHITECTURE arc OF MAQUINA_DE_ESTADOS IS
	TYPE ESTADO IS ( REALIZAR_AMOSTRAGEM, AGUARDAR );
	SIGNAL shift_reg :STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL state : ESTADO := REALIZAR_AMOSTRAGEM;
BEGIN

PROCESS(clk) IS
	VARIABLE cont: INTEGER := 0 ;
BEGIN
	IF RISING_EDGE(clk) THEN
		CASE state IS
			WHEN REALIZAR_AMOSTRAGEM =>
				shift_reg(7) <= botao;
				shift_reg(6 DOWNTO 0) <= shift_reg(7 DOWNTO 1);
				state <= AGUARDAR;
			WHEN AGUARDAR =>
		--	3333333
				IF cont < 333333 THEN
					cont:= cont + 1;
				ELSIF cont = 333333 THEN
					cont:=0;
					state <= REALIZAR_AMOSTRAGEM;
				END IF;
		END CASE;
	
		IF shift_reg = "11111111" THEN
			saida<= '1';
		ELSIF shift_reg = "00000000" THEN
			saida<='0';
		ELSE
			saida<=saida;
		END IF;
	END IF;
END PROCESS;

END ARCHITECTURE;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE pacotin IS

COMPONENT  MAQUINA_DE_ESTADOS IS
	PORT (botao,clk: IN  STD_LOGIC;
          saida:BUFFER STD_LOGIC);
END COMPONENT;

END PACKAGE;