LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY DIVISOR_DE_FREQUENCIA IS
	GENERIC(cont:INTEGER:=10);
	PORT(clk66:IN STD_LOGIC;
		 clk_dividido:BUFFER STD_LOGIC);
END ENTITY;

ARCHITECTURE arc OF DIVISOR_DE_FREQUENCIA IS
BEGIN
	PROCESS(clk66) IS
		VARIABLE c:INTEGER := 0;
	BEGIN
		IF RISING_EDGE(clk66) THEN
			c := c + 1;
			IF c = cont THEN
				c := 0;
				clk_dividido<=NOT clk_dividido;
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE;