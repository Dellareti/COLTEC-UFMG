--LIBRARY IEEE;
--USE IEEE.STD_LOGIC_1164.ALL;
--USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--USE IEEE.NUMERIC_STD.ALL;
--USE IEEE.STD_LOGIC_ARITH.ALL;
--USE WORK.COMPONENTES.ALL;
--
--ENTITY TOP_ENTITY IS
--
--END ENTITY;
--
--ARCHITECTURE top_design OF TOP_ENTITY IS
--BEGIN
--
--END ARCHITECTURE;